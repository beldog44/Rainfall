b0VIM 7.3      q�XT�T5  t-kamano                                softbank126017073004.bbtec.net          ~t-kamano/test_company/tutorial/tutorial/spiders/webspider.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ad  O
  �
             �  �  �  �  �  ]  \  6    �  �  k  F    �  �  �  �  0    �  `  5  +      �  �  �  F     �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          yield article        #article['name'] = response.css("td.data_0_0").extract_first()               yield article        #article['name'] = response.css("td.data_0_0").extract_first()        # article['time']  = response.css("td.white-space:nowrap").extract_first()        article['time']  = response.xpath('//td/text()').extract()        article = WebItem()     def parse(self, response):          print ('end')     else:         #d1 + datetime.timedelta(days = 1) 	start_urls = ['http://www.data.jma.go.jp/obd/stats/etrn/view/10min_s1.php?prec_no=62&block_no=47772&year=2017&month=03&day={0}&view=a4'.format(dd1)] 	dd1 = (d1.day)         d1 + datetime.timedelta(days = 1)         #dd1 = (d1.day)                #繰り返す度に日付を更新するため         print ('start')     if d1 <= d2:     #td = datetime.timedelta(days=1)  #for文で回るようにする     #print (d1)     d2 = date(2017, 3, 31)                #調査最終年月日     #d = datetime.date(20:16, 6, 27)     dd1 = (d1.day)                        #調査日付のみ     d1 = date(2017, 3, 29)                #調査年月日     allowed_domains = ["http://www.data.jma.go.jp/"]     name = "webspiderSpider" class WebSpiderSpider(scrapy.Spider):  from scrapy.linkextractors import LinkExtractor from tutorial.items import WebItem from datetime import date import datetime import scrapy # -*- coding: utf-8 -*- 